`include "abs.vh"
`include "log2.vh"
